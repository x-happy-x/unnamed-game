[MENU PAUSE] - Элементы меню паузы
ПРОДОЛЖИТЬ
НАЧАТЬ СНАЧАЛО
ПРОПУСТИТЬ УРОВЕНЬ
ОТЧЁТ ОБ ОШИБКЕ
ГЛАВНОЕ МЕНЮ

[MENU END] - Элементы меню в конце игры
ДАЛЕЕ
НАЧАТЬ СНАЧАЛО
ОТЧЁТ ОБ ОШИБКЕ
ГЛАВНОЕ МЕНЮ

[USE HELP] - Когда использовал подсказку
[MusicLevel] Теперь вы можете слушать песню полностью
[Aesthetics] Открыта дополнительная картинка

[USE TICKET] - Когда использовал пропуск
[MusicLevel] Хммммм так не честно
[Aesthetics] Хммммм так не честно

[USED HELP] - Когда уже использовал подсказку
Ну чего тебе?_Ты уже использовал её
Вы уже использовали её
Вы уже воспользовались подсказкой

[ERROR] - Надпись при неправильном ответе
Ты по своему прав, а по-моему нет
Не верно, дурак :)
Неправильно, бугага

[ERROR COUNT] - Когда несколько ошибок отнимают жизнь
[FIRST]Помни! {0} - минус жизнь
[FIRST]Не забудь, что {0} отнимут жизнь!
[OTHER]Ещё {1} и мне наскучит
[END]{2} хорошо, но и {3} неплохо

[WIN] - Надпись при правильном ответе (от 1 до 5 степень правильности)
[5]Идеально
[4]Отличненько
[3]Ух ты ж пух ты
[2]Нууу ладно, верно
[1]Верно, но всё равно дурак :)
[0]Если ты видишь это, то ты__ что-то скрываешь -_-

[WIN HELP] - Надпись при правильном ответе с использованием подсказки
Ай яй яй, с подсказками только и можешь
Ах ты ж жулик
Ну так кто угодно сможет
Правильно... P.S. но я знаю что ты жулик :)

[NO TICKET] - Когда нет пропусков
Ууупс у вас закончились пропуски
Хихихи, а их у вас нет
Ну нет их, что ты хочешь?

[NO HELP] - Когда нет подсказок
Я бы отдал, но где их взять
А не жирно ли будет?
Ага, раскатал губу
Вы не расстраивайтесь,__но они закончились :(

[NO LIVE] - Когда нет жизней
Я бы отдал, но где их взять
А не жирно ли будет?
Ага, раскатал губу
Вы не расстраивайтесь,__но они закончились :(

[NO LEVEL] - Когда нет следующего уровня
Уууууууууупс, а его нет

[NO TEXT] - Когда не ввели текст
Вы не ввели ничего
Вы не ввели текст

[click for retry] - Для переподключения
Нажмите на экран чтобы попробовать снова